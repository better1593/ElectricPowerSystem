* netlist generated with vector fitting poles and residues

.subckt total_network node_1 node_2 node_3 node_ref
X_11 node_1 node_ref yp11
X_12 node_1 node_2 yp12
X_13 node_1 node_3 yp13
X_22 node_2 node_ref yp22
X_23 node_2 node_3 yp23
X_33 node_3 node_ref yp33
.ends


* Y'11
.subckt yp11 node_1 node_ref
* Branch 0
Rabr0 node_1 netRa0 104.85192466442048
Lbr0 netRa0 netL0 0.03603571280837059
Rbbr0 netL0 node_ref 66538.29858456686
Cbr0 netL0 node_ref 2.221486955304943e-08

* Branch 1
Rabr1 node_1 netRa1 23.97092422447678
Lbr1 netRa1 netL1 0.01655505783855915
Rbbr1 netL1 node_ref 24314.77955789861
Cbr1 netL1 node_ref 3.998093983020541e-08

* Branch 2
Rabr2 node_1 netRa2 -80.53191078383787
Lbr2 netRa2 netL2 0.0430884063243866
Rbbr2 netL2 node_ref -28481.82621995759
Cbr2 netL2 node_ref 1.514039473324074e-08

* Branch 3
Rabr3 node_1 netRa3 284.7911106620841
Lbr3 netRa3 netL3 0.03451797738671303
Rbbr3 netL3 node_ref 266153.1416134351
Cbr3 netL3 node_ref 2.463498888694679e-09

* Branch 4
Rabr4 node_1 netRa4 51.35181677247574
Lbr4 netRa4 netL4 0.01661824993789196
Rbbr4 netL4 node_ref 98263.51501565707
Cbr4 netL4 node_ref 4.404482496919189e-09

* Branch 5
Rabr5 node_1 netRa5 -133.93483142158516
Lbr5 netRa5 netL5 0.04242291674017906
Rbbr5 netL5 node_ref -149592.78834168628
Cbr5 netL5 node_ref 1.7061983924393958e-09

* Branch 6
Rabr6 node_1 netRa6 476.9334390075544
Lbr6 netRa6 netL6 0.033604610711336136
Rbbr6 netL6 node_ref 359310.375907067
Cbr6 netL6 node_ref 8.924682559742155e-10

* Branch 7
Rabr7 node_1 netRa7 110.96724584478416
Lbr7 netRa7 netL7 0.01580631360411644
Rbbr7 netL7 node_ref 102498.09162027646
Cbr7 netL7 node_ref 1.662917287657302e-09

* Branch 8
Rabr8 node_1 netRa8 -596.6858836538272
Lbr8 netRa8 netL8 0.04729977250099182
Rbbr8 netL8 node_ref -134389.70192382723
Cbr8 netL8 node_ref 5.48686756683558e-10

* Branch 9
Rabr9 node_1 netRa9 577.5568832916686
Lbr9 netRa9 netL9 0.03249189257621765
Rbbr9 netL9 node_ref 855330.5591527633
Cbr9 netL9 node_ref 4.6460874302326943e-10

* Branch 10
Rabr10 node_1 netRa10 61.07271315221466
Lbr10 netRa10 netL10 0.015984030440449715
Rbbr10 netL10 node_ref 507457.2168351258
Cbr10 netL10 node_ref 8.389822207433891e-10

* Branch 11
Rabr11 node_1 netRa11 111.29626450858697
Lbr11 netRa11 netL11 0.04468223825097084
Rbbr11 netL11 node_ref 2499265.822551149
Cbr11 netL11 node_ref 2.97449223919291e-10

* Branch 12
Rabr12 node_1 netRa12 609.246825849404
Lbr12 netRa12 netL12 0.031282681971788406
Rbbr12 netL12 node_ref 61028624.02375445
Cbr12 netL12 node_ref 2.8909752985160475e-10

* Branch 13
Rabr13 node_1 netRa13 103.61963736973688
Lbr13 netRa13 netL13 0.01568642258644104
Rbbr13 netL13 node_ref 406239.2500308092
Cbr13 netL13 node_ref 5.167552336953745e-10

* Branch 14
Rabr14 node_1 netRa14 51.50012020780365
Lbr14 netRa14 netL14 0.04599593207240105
Rbbr14 netL14 node_ref -40290937.88077229
Cbr14 netL14 node_ref 1.747381220613374e-10

* Branch 15
Rabr15 node_1 netRa15 466.09937405983766
Lbr15 netRa15 netL15 0.030966438353061676
Rbbr15 netL15 node_ref -653521.8212227856
Cbr15 netL15 node_ref 1.940565573658753e-10

* Branch 16
Rabr16 node_1 netRa16 36.20229772498286
Lbr16 netRa16 netL16 0.015594634227454662
Rbbr16 netL16 node_ref 19957307.02570276
Cbr16 netL16 node_ref 3.4782298578574673e-10

* Branch 17
Rabr17 node_1 netRa17 802.21013722832
Lbr17 netRa17 netL17 0.04518767446279526
Rbbr17 netL17 node_ref 514865.8899008287
Cbr17 netL17 node_ref 1.1883822778727674e-10

* Branch 18
Rabr18 node_1 netRa18 -772.8739795137145
Lbr18 netRa18 netL18 0.03216779604554176
Rbbr18 netL18 node_ref -152609.6954652635
Cbr18 netL18 node_ref 1.3192331402624544e-10

* Branch 19
Rabr19 node_1 netRa19 -106.60960160781026
Lbr19 netRa19 netL19 0.015438985079526901
Rbbr19 netL19 node_ref -422236.21560827084
Cbr19 netL19 node_ref 2.5131929904167295e-10

* Branch 20
Rabr20 node_1 netRa20 1910.1162684640065
Lbr20 netRa20 netL20 0.04415206238627434
Rbbr20 netL20 node_ref 277026.0023609452
Cbr20 netL20 node_ref 8.659131497775039e-11

* Branch 21
Rabr21 node_1 netRa21 -6414.511672807723
Lbr21 netRa21 netL21 0.03976304829120636
Rbbr21 netL21 node_ref -73293.8166760016
Cbr21 netL21 node_ref 7.289610629705023e-11

* Branch 22
Rabr22 node_1 netRa22 -321.9703869967046
Lbr22 netRa22 netL22 0.015935653820633888
Rbbr22 netL22 node_ref -238240.7991738014
Cbr22 netL22 node_ref 1.8259449141475423e-10

* Branch 23
Rabr23 node_1 netRa23 1659.6221779954433
Lbr23 netRa23 netL23 0.04173152521252632
Rbbr23 netL23 node_ref 381421.1098806523
Cbr23 netL23 node_ref 6.89703224296523e-11

* Branch 24
Rabr24 node_1 netRa24 572.7548833898331
Lbr24 netRa24 netL24 0.0010093661257997155
Rbbr24 netL24 node_ref 2018.6334125094236
Cbr24 netL24 node_ref 1.2626807262004068e-09

.ends


* Y'12
.subckt yp12 node_1 node_2
* Branch 0
Rabr0 node_1 netRa0 103.64695364114418
Lbr0 netRa0 netL0 0.04196883738040924
Rbbr0 netL0 node_2 221452.70573922823
Cbr0 netL0 node_2 1.909552166209675e-08

* Branch 1
Rabr1 node_1 netRa1 -969.3807679012154
Lbr1 netRa1 netL1 -0.11989299952983856
Rbbr1 netL1 node_2 -24574.552164284978
Cbr1 netL1 node_2 -5.3081076050630615e-09

* Branch 2
Rabr2 node_1 netRa2 21.32685628231911
Lbr2 netRa2 netL2 -0.026652611792087555
Rbbr2 netL2 node_2 32608.636317867215
Cbr2 netL2 node_2 -2.4530333180030658e-08

* Branch 3
Rabr3 node_1 netRa3 189.82817231301047
Lbr3 netRa3 netL3 0.04020218551158905
Rbbr3 netL3 node_2 -235528.94481300714
Cbr3 netL3 node_2 2.1191556257871717e-09

* Branch 4
Rabr4 node_1 netRa4 -16864.19599551901
Lbr4 netRa4 netL4 -0.32824334502220154
Rbbr4 netL4 node_2 -105448.97195509999
Cbr4 netL4 node_2 -1.8742522533146923e-10

* Branch 5
Rabr5 node_1 netRa5 31.43070600883335
Lbr5 netRa5 netL5 -0.023179588839411736
Rbbr5 netL5 node_2 151181.71660450907
Cbr5 netL5 node_2 -3.1248059747703855e-09

* Branch 6
Rabr6 node_1 netRa6 301.0445579573902
Lbr6 netRa6 netL6 0.03967059403657913
Rbbr6 netL6 node_2 -378700.5870635287
Cbr6 netL6 node_2 7.576085705108785e-10

* Branch 7
Rabr7 node_1 netRa7 -70936.37585270617
Lbr7 netRa7 netL7 -1.1382427215576172
Rbbr7 netL7 node_2 -778136.8768196767
Cbr7 netL7 node_2 -2.1009870438296982e-11

* Branch 8
Rabr8 node_1 netRa8 -90.7655265056904
Lbr8 netRa8 netL8 -0.021878574043512344
Rbbr8 netL8 node_2 -262197.0611439022
Cbr8 netL8 node_2 -1.1910958259899833e-09

* Branch 9
Rabr9 node_1 netRa9 267.7821616617235
Lbr9 netRa9 netL9 0.0395892858505249
Rbbr9 netL9 node_2 -308234.02262650826
Cbr9 netL9 node_2 3.8190494017008186e-10

* Branch 10
Rabr10 node_1 netRa10 -875921.8318175554
Lbr10 netRa10 netL10 -2.2611193656921387
Rbbr10 netL10 node_2 -1312783.2871040606
Cbr10 netL10 node_2 -1.9738699346550394e-12

* Branch 11
Rabr11 node_1 netRa11 -89.74124836200558
Lbr11 netRa11 netL11 -0.021566342562437057
Rbbr11 netL11 node_2 -538174.5245200521
Cbr11 netL11 node_2 -6.161950528235442e-10

* Branch 12
Rabr12 node_1 netRa12 344.18174318454936
Lbr12 netRa12 netL12 0.039859481155872345
Rbbr12 netL12 node_2 -408351.6100822344
Cbr12 netL12 node_2 2.27084194236278e-10

* Branch 13
Rabr13 node_1 netRa13 -51622.06527723762
Lbr13 netRa13 netL13 -0.7625031471252441
Rbbr13 netL13 node_2 -1479558.9302112667
Cbr13 netL13 node_2 -1.0262536387940108e-11

* Branch 14
Rabr14 node_1 netRa14 -231.0067361960215
Lbr14 netRa14 netL14 -0.021792376413941383
Rbbr14 netL14 node_2 -290575.9997900529
Cbr14 netL14 node_2 -3.685161419102135e-10

* Branch 15
Rabr15 node_1 netRa15 403.1893622444254
Lbr15 netRa15 netL15 0.0412612222135067
Rbbr15 netL15 node_2 -521513.45799074415
Cbr15 netL15 node_2 1.4564762116081024e-10

* Branch 16
Rabr16 node_1 netRa16 -27884.980101315392
Lbr16 netRa16 netL16 -0.7510207891464233
Rbbr16 netL16 node_2 -3989252.9968086057
Cbr16 netL16 node_2 -7.171928288131466e-12

* Branch 17
Rabr17 node_1 netRa17 -295.3293497135498
Lbr17 netRa17 netL17 -0.02166745997965336
Rbbr17 netL17 node_2 -329943.8932252704
Cbr17 netL17 node_2 -2.4800273993421895e-10

* Branch 18
Rabr18 node_1 netRa18 321.47840202832754
Lbr18 netRa18 netL18 0.04442785680294037
Rbbr18 netL18 node_2 -565529.2190635762
Cbr18 netL18 node_2 9.605927537903679e-11

* Branch 19
Rabr19 node_1 netRa19 318802.5063019276
Lbr19 netRa19 netL19 -1.2547166347503662
Rbbr19 netL19 node_2 1578690.1670666512
Cbr19 netL19 node_2 -2.468559311786439e-12

* Branch 20
Rabr20 node_1 netRa20 -374.07217887182776
Lbr20 netRa20 netL20 -0.021255237981677055
Rbbr20 netL20 node_2 -344928.26773976313
Cbr20 netL20 node_2 -1.809226594200938e-10

* Branch 21
Rabr21 node_1 netRa21 13.386181570598286
Lbr21 netRa21 netL21 0.05302750691771507
Rbbr21 netL21 node_2 -652176.419323957
Cbr21 netL21 node_2 5.990558386475362e-11

* Branch 22
Rabr22 node_1 netRa22 2965272.522889833
Lbr22 netRa22 netL22 1.6699694395065308
Rbbr22 netL22 node_2 3288559.9434428643
Cbr22 netL22 node_2 1.7152184314631018e-13

* Branch 23
Rabr23 node_1 netRa23 -252.2272019300616
Lbr23 netRa23 netL23 -0.02032398246228695
Rbbr23 netL23 node_2 -660125.7744863468
Cbr23 netL23 node_2 -1.4218229993436607e-10

* Branch 24
Rabr24 node_1 netRa24 -1188152.3894957248
Lbr24 netRa24 netL24 0.07660263776779175
Rbbr24 netL24 node_2 -1190896.8406592226
Cbr24 netL24 node_2 5.353301980876685e-14

.ends


* Y'13
.subckt yp13 node_1 node_3
* Branch 0
Rabr0 node_1 netRa0 82.60251111840002
Lbr0 netRa0 netL0 0.03599238023161888
Rbbr0 netL0 node_3 725765.8418849265
Cbr0 netL0 node_3 2.22741803708322e-08

* Branch 1
Rabr1 node_1 netRa1 -45.42836309481833
Lbr1 netRa1 netL1 -0.01936163380742073
Rbbr1 netL1 node_3 -15210.411108099055
Cbr1 netL1 node_3 -3.411701088475873e-08

* Branch 2
Rabr2 node_1 netRa2 652.6747369170425
Lbr2 netRa2 netL2 0.08113505691289902
Rbbr2 netL2 node_3 16982.89749181778
Cbr2 netL2 node_3 7.753523052921687e-09

* Branch 3
Rabr3 node_1 netRa3 150.23065429235348
Lbr3 netRa3 netL3 0.034838609397411346
Rbbr3 netL3 node_3 -169444.04515916665
Cbr3 netL3 node_3 2.445607366858725e-09

* Branch 4
Rabr4 node_1 netRa4 -28.95151191368231
Lbr4 netRa4 netL4 -0.017462877556681633
Rbbr4 netL4 node_3 -271514.0878592472
Cbr4 netL4 node_3 -4.1931950869178334e-09

* Branch 5
Rabr5 node_1 netRa5 147.45222280403746
Lbr5 netRa5 netL5 0.056068502366542816
Rbbr5 netL5 node_3 414226.05642333196
Cbr5 netL5 node_3 1.2916519533276192e-09

* Branch 6
Rabr6 node_1 netRa6 252.9707715581498
Lbr6 netRa6 netL6 0.03457454591989517
Rbbr6 netL6 node_3 -306156.76400491886
Cbr6 netL6 node_3 8.693019960198051e-10

* Branch 7
Rabr7 node_1 netRa7 -111.17191014225288
Lbr7 netRa7 netL7 -0.01582586020231247
Rbbr7 netL7 node_3 -102550.50578806213
Cbr7 netL7 node_3 -1.6608610551419188e-09

* Branch 8
Rabr8 node_1 netRa8 503.1464917457077
Lbr8 netRa8 netL8 0.04228358343243599
Rbbr8 netL8 node_3 148595.29919874266
Cbr8 netL8 node_3 6.144283987476824e-10

* Branch 9
Rabr9 node_1 netRa9 256.68513047311586
Lbr9 netRa9 netL9 0.034447863698005676
Rbbr9 netL9 node_3 -291814.22885175416
Cbr9 netL9 node_3 4.3890982057571203e-10

* Branch 10
Rabr10 node_1 netRa10 -101.62279376439128
Lbr10 netRa10 netL10 -0.015954019501805305
Rbbr10 netL10 node_3 -242979.67557093364
Cbr10 netL10 node_3 -8.403100457010613e-10

* Branch 11
Rabr11 node_1 netRa11 285.7934562160289
Lbr11 netRa11 netL11 0.04341292008757591
Rbbr11 netL11 node_3 600982.5751874038
Cbr11 netL11 node_3 3.060141862468441e-10

* Branch 12
Rabr12 node_1 netRa12 330.80123914888225
Lbr12 netRa12 netL12 0.034602291882038116
Rbbr12 netL12 node_3 -387757.0971996305
Cbr12 netL12 node_3 2.6158823340242216e-10

* Branch 13
Rabr13 node_1 netRa13 -187.48463714004808
Lbr13 netRa13 netL13 -0.015834981575608253
Rbbr13 netL13 node_3 -195528.7216743811
Cbr13 netL13 node_3 -5.11546820436068e-10

* Branch 14
Rabr14 node_1 netRa14 618.3622401339288
Lbr14 netRa14 netL14 0.04266473278403282
Rbbr14 netL14 node_3 401801.8023594529
Cbr14 netL14 node_3 1.8809127066015914e-10

* Branch 15
Rabr15 node_1 netRa15 456.5409113898496
Lbr15 netRa15 netL15 0.03545800969004631
Rbbr15 netL15 node_3 -586418.9436278228
Cbr15 netL15 node_3 1.6948586570047103e-10

* Branch 16
Rabr16 node_1 netRa16 -162.8162841423711
Lbr16 netRa16 netL16 -0.015819786116480827
Rbbr16 netL16 node_3 -359582.9383093282
Cbr16 netL16 node_3 -3.427180867489614e-10

* Branch 17
Rabr17 node_1 netRa17 346.04744279033525
Lbr17 netRa17 netL17 0.04291946068406105
Rbbr17 netL17 node_3 1199702.346775848
Cbr17 netL17 node_3 1.252777089416227e-10

* Branch 18
Rabr18 node_1 netRa18 501.8926486702683
Lbr18 netRa18 netL18 0.037774261087179184
Rbbr18 netL18 node_3 -716177.2066677687
Cbr18 netL18 node_3 1.1299419718699155e-10

* Branch 19
Rabr19 node_1 netRa19 -47.90607861889786
Lbr19 netRa19 netL19 -0.015585231594741344
Rbbr19 netL19 node_3 -7230376.088335858
Cbr19 netL19 node_3 -2.490222272622208e-10

* Branch 20
Rabr20 node_1 netRa20 -318.5964759302626
Lbr20 netRa20 netL20 0.04222247004508972
Rbbr20 netL20 node_3 -1202852.1001239384
Cbr20 netL20 node_3 9.115311605462798e-11

* Branch 21
Rabr21 node_1 netRa21 -150.80875221681072
Lbr21 netRa21 netL21 0.044867683202028275
Rbbr21 netL21 node_3 -483712.60104352544
Cbr21 netL21 node_3 7.077673274388957e-11

* Branch 22
Rabr22 node_1 netRa22 321.34791391703254
Lbr22 netRa22 netL22 -0.015583254396915436
Rbbr22 netL22 node_3 228834.02506765444
Cbr22 netL22 node_3 -1.8671383301141504e-10

* Branch 23
Rabr23 node_1 netRa23 -841.6983725179946
Lbr23 netRa23 netL23 0.04325864836573601
Rbbr23 netL23 node_3 -706256.3454829996
Cbr23 netL23 node_3 6.674665555347314e-11

* Branch 24
Rabr24 node_1 netRa24 -25841.266547787258
Lbr24 netRa24 netL24 0.01300709880888462
Rbbr24 netL24 node_3 -29222.643066460045
Cbr24 netL24 node_3 1.582929148560598e-11

.ends


* Y'22
.subckt yp22 node_2 node_ref
* Branch 0
Rabr0 node_2 netRa0 201.0954228197926
Lbr0 netRa0 netL0 0.04851918667554855
Rbbr0 netL0 node_ref 31858.37775142082
Cbr0 netL0 node_ref 1.6420946209881034e-08

* Branch 1
Rabr1 node_2 netRa1 149.98934173169351
Lbr1 netRa1 netL1 0.05436384677886963
Rbbr1 netL1 node_ref 35220.01332292542
Cbr1 netL1 node_ref 1.2135240185470451e-08

* Branch 2
Rabr2 node_2 netRa2 -1.7905573401330008
Lbr2 netRa2 netL2 0.012692018412053585
Rbbr2 netL2 node_ref -32824.64860955008
Cbr2 netL2 node_ref 5.154338336962283e-08

* Branch 3
Rabr3 node_2 netRa3 628.6170971647808
Lbr3 netRa3 netL3 0.04563424363732338
Rbbr3 netL3 node_ref 76670.6237078725
Cbr3 netL3 node_ref 1.8501049933810875e-09

* Branch 4
Rabr4 node_2 netRa4 6457.487313008619
Lbr4 netRa4 netL4 0.15647096931934357
Rbbr4 netL4 node_ref 59226.47335957143
Cbr4 netL4 node_ref 4.1700024595623006e-10

* Branch 5
Rabr5 node_2 netRa5 -28.07835474176541
Lbr5 netRa5 netL5 0.011055068112909794
Rbbr5 netL5 node_ref -46259.571467802416
Cbr5 netL5 node_ref 6.5492867831288714e-09

* Branch 6
Rabr6 node_2 netRa6 1081.3756026003934
Lbr6 netRa6 netL6 0.043877094984054565
Rbbr6 netL6 node_ref 108738.16253090023
Cbr6 netL6 node_ref 6.776260006131186e-10

* Branch 7
Rabr7 node_2 netRa7 45433.616048368065
Lbr7 netRa7 netL7 0.8822208046913147
Rbbr7 netL7 node_ref 711386.4888748797
Cbr7 netL7 node_ref 2.7921080492240425e-11

* Branch 8
Rabr8 node_2 netRa8 -1.3356220485036592
Lbr8 netRa8 netL8 0.010387214832007885
Rbbr8 netL8 node_ref -370606.47449026123
Cbr8 netL8 node_ref 2.5096629215702196e-09

* Branch 9
Rabr9 node_2 netRa9 1334.669825350862
Lbr9 netRa9 netL9 0.04160981625318527
Rbbr9 netL9 node_ref 165127.947416389
Cbr9 netL9 node_ref 3.601102432215579e-10

* Branch 10
Rabr10 node_2 netRa10 267736.7089706317
Lbr10 netRa10 netL10 2.2658591270446777
Rbbr10 netL10 node_ref 1715544.810172989
Cbr10 netL10 node_ref 4.995366584820152e-12

* Branch 11
Rabr11 node_2 netRa11 4.000894428396884
Lbr11 netRa11 netL11 0.010277559980750084
Rbbr11 netL11 node_ref -1022290.0533532389
Cbr11 netL11 node_ref 1.2932391437738751e-09

* Branch 12
Rabr12 node_2 netRa12 1434.1316607407907
Lbr12 netRa12 netL12 0.03935174643993378
Rbbr12 netL12 node_ref 257011.62687929862
Cbr12 netL12 node_ref 2.285380525415859e-10

* Branch 13
Rabr13 node_2 netRa13 -46935.30505781771
Lbr13 netRa13 netL13 0.4724588096141815
Rbbr13 netL13 node_ref -622811.7180280111
Cbr13 netL13 node_ref 1.5868219063779582e-11

* Branch 14
Rabr14 node_2 netRa14 45.67890005129542
Lbr14 netRa14 netL14 0.01038623508065939
Rbbr14 netL14 node_ref 412078.23142775433
Cbr14 netL14 node_ref 7.737492157703496e-10

* Branch 15
Rabr15 node_2 netRa15 1311.447069300252
Lbr15 netRa15 netL15 0.03808590769767761
Rbbr15 netL15 node_ref 552970.4622200334
Cbr15 netL15 node_ref 1.572948010867124e-10

* Branch 16
Rabr16 node_2 netRa16 -72708.11605479202
Lbr16 netRa16 netL16 0.4147893488407135
Rbbr16 netL16 node_ref -503608.1687268674
Cbr16 netL16 node_ref 1.1188978536366796e-11

* Branch 17
Rabr17 node_2 netRa17 71.34261563744124
Lbr17 netRa17 netL17 0.010349337942898273
Rbbr17 netL17 node_ref 350936.6704375168
Cbr17 netL17 node_ref 5.195800806323321e-10

* Branch 18
Rabr18 node_2 netRa18 -171.0374227991533
Lbr18 netRa18 netL18 0.03877369314432144
Rbbr18 netL18 node_ref -302633.2903437948
Cbr18 netL18 node_ref 1.0994239127958196e-10

* Branch 19
Rabr19 node_2 netRa19 -388609.12230937975
Lbr19 netRa19 netL19 0.6824701428413391
Rbbr19 netL19 node_ref -696065.495575837
Cbr19 netL19 node_ref 2.5119098806103e-12

* Branch 20
Rabr20 node_2 netRa20 99.84737804738222
Lbr20 netRa20 netL20 0.01016842108219862
Rbbr20 netL20 node_ref 320472.3780755693
Cbr20 netL20 node_ref 3.7847861700717583e-10

* Branch 21
Rabr21 node_2 netRa21 -7598.560315614798
Lbr21 netRa21 netL21 0.047556985169649124
Rbbr21 netL21 node_ref -88250.62623027405
Cbr21 netL21 node_ref 6.104399586359392e-11

* Branch 22
Rabr22 node_2 netRa22 -265724.7360347152
Lbr22 netRa22 netL22 -0.47269490361213684
Rbbr22 netL22 node_ref -555753.1507241023
Cbr22 netL22 node_ref -3.2167891313152335e-12

* Branch 23
Rabr23 node_2 netRa23 24.907236864556335
Lbr23 netRa23 netL23 0.009861026890575886
Rbbr23 netL23 node_ref 4430834.964342797
Cbr23 netL23 node_ref 2.9315393799561067e-10

* Branch 24
Rabr24 node_2 netRa24 652.1448658077649
Lbr24 netRa24 netL24 0.0010242159478366375
Rbbr24 netL24 node_ref 1899.0836227172304
Cbr24 netL24 node_ref 1.1407157692238187e-09

.ends


* Y'23
.subckt yp23 node_2 node_3
* Branch 0
Rabr0 node_2 netRa0 103.64695364114418
Lbr0 netRa0 netL0 0.04196883738040924
Rbbr0 netL0 node_3 221452.70573922823
Cbr0 netL0 node_3 1.909552166209675e-08

* Branch 1
Rabr1 node_2 netRa1 -969.3807679012154
Lbr1 netRa1 netL1 -0.11989299952983856
Rbbr1 netL1 node_3 -24574.552164284978
Cbr1 netL1 node_3 -5.3081076050630615e-09

* Branch 2
Rabr2 node_2 netRa2 21.32685628231911
Lbr2 netRa2 netL2 -0.026652611792087555
Rbbr2 netL2 node_3 32608.636317867215
Cbr2 netL2 node_3 -2.4530333180030658e-08

* Branch 3
Rabr3 node_2 netRa3 189.82817231301047
Lbr3 netRa3 netL3 0.04020218551158905
Rbbr3 netL3 node_3 -235528.94481300714
Cbr3 netL3 node_3 2.1191556257871717e-09

* Branch 4
Rabr4 node_2 netRa4 -16864.19599551901
Lbr4 netRa4 netL4 -0.32824334502220154
Rbbr4 netL4 node_3 -105448.97195509999
Cbr4 netL4 node_3 -1.8742522533146923e-10

* Branch 5
Rabr5 node_2 netRa5 31.43070600883335
Lbr5 netRa5 netL5 -0.023179588839411736
Rbbr5 netL5 node_3 151181.71660450907
Cbr5 netL5 node_3 -3.1248059747703855e-09

* Branch 6
Rabr6 node_2 netRa6 301.0445579573902
Lbr6 netRa6 netL6 0.03967059403657913
Rbbr6 netL6 node_3 -378700.5870635287
Cbr6 netL6 node_3 7.576085705108785e-10

* Branch 7
Rabr7 node_2 netRa7 -70936.37585270617
Lbr7 netRa7 netL7 -1.1382427215576172
Rbbr7 netL7 node_3 -778136.8768196767
Cbr7 netL7 node_3 -2.1009870438296982e-11

* Branch 8
Rabr8 node_2 netRa8 -90.7655265056904
Lbr8 netRa8 netL8 -0.021878574043512344
Rbbr8 netL8 node_3 -262197.0611439022
Cbr8 netL8 node_3 -1.1910958259899833e-09

* Branch 9
Rabr9 node_2 netRa9 267.7821616617235
Lbr9 netRa9 netL9 0.0395892858505249
Rbbr9 netL9 node_3 -308234.02262650826
Cbr9 netL9 node_3 3.8190494017008186e-10

* Branch 10
Rabr10 node_2 netRa10 -875921.8318175554
Lbr10 netRa10 netL10 -2.2611193656921387
Rbbr10 netL10 node_3 -1312783.2871040606
Cbr10 netL10 node_3 -1.9738699346550394e-12

* Branch 11
Rabr11 node_2 netRa11 -89.74124836200558
Lbr11 netRa11 netL11 -0.021566342562437057
Rbbr11 netL11 node_3 -538174.5245200521
Cbr11 netL11 node_3 -6.161950528235442e-10

* Branch 12
Rabr12 node_2 netRa12 344.18174318454936
Lbr12 netRa12 netL12 0.039859481155872345
Rbbr12 netL12 node_3 -408351.6100822344
Cbr12 netL12 node_3 2.27084194236278e-10

* Branch 13
Rabr13 node_2 netRa13 -51622.06527723762
Lbr13 netRa13 netL13 -0.7625031471252441
Rbbr13 netL13 node_3 -1479558.9302112667
Cbr13 netL13 node_3 -1.0262536387940108e-11

* Branch 14
Rabr14 node_2 netRa14 -231.0067361960215
Lbr14 netRa14 netL14 -0.021792376413941383
Rbbr14 netL14 node_3 -290575.9997900529
Cbr14 netL14 node_3 -3.685161419102135e-10

* Branch 15
Rabr15 node_2 netRa15 403.1893622444254
Lbr15 netRa15 netL15 0.0412612222135067
Rbbr15 netL15 node_3 -521513.45799074415
Cbr15 netL15 node_3 1.4564762116081024e-10

* Branch 16
Rabr16 node_2 netRa16 -27884.980101315392
Lbr16 netRa16 netL16 -0.7510207891464233
Rbbr16 netL16 node_3 -3989252.9968086057
Cbr16 netL16 node_3 -7.171928288131466e-12

* Branch 17
Rabr17 node_2 netRa17 -295.3293497135498
Lbr17 netRa17 netL17 -0.02166745997965336
Rbbr17 netL17 node_3 -329943.8932252704
Cbr17 netL17 node_3 -2.4800273993421895e-10

* Branch 18
Rabr18 node_2 netRa18 321.47840202832754
Lbr18 netRa18 netL18 0.04442785680294037
Rbbr18 netL18 node_3 -565529.2190635762
Cbr18 netL18 node_3 9.605927537903679e-11

* Branch 19
Rabr19 node_2 netRa19 318802.5063019276
Lbr19 netRa19 netL19 -1.2547166347503662
Rbbr19 netL19 node_3 1578690.1670666512
Cbr19 netL19 node_3 -2.468559311786439e-12

* Branch 20
Rabr20 node_2 netRa20 -374.07217887182776
Lbr20 netRa20 netL20 -0.021255237981677055
Rbbr20 netL20 node_3 -344928.26773976313
Cbr20 netL20 node_3 -1.809226594200938e-10

* Branch 21
Rabr21 node_2 netRa21 13.386181570598286
Lbr21 netRa21 netL21 0.05302750691771507
Rbbr21 netL21 node_3 -652176.419323957
Cbr21 netL21 node_3 5.990558386475362e-11

* Branch 22
Rabr22 node_2 netRa22 2965272.522889833
Lbr22 netRa22 netL22 1.6699694395065308
Rbbr22 netL22 node_3 3288559.9434428643
Cbr22 netL22 node_3 1.7152184314631018e-13

* Branch 23
Rabr23 node_2 netRa23 -252.2272019300616
Lbr23 netRa23 netL23 -0.02032398246228695
Rbbr23 netL23 node_3 -660125.7744863468
Cbr23 netL23 node_3 -1.4218229993436607e-10

* Branch 24
Rabr24 node_2 netRa24 -1188152.3894957248
Lbr24 netRa24 netL24 0.07660263776779175
Rbbr24 netL24 node_3 -1190896.8406592226
Cbr24 netL24 node_3 5.353301980876685e-14

.ends


* Y'33
.subckt yp33 node_3 node_ref
* Branch 0
Rabr0 node_3 netRa0 104.85192466442048
Lbr0 netRa0 netL0 0.03603571280837059
Rbbr0 netL0 node_ref 66538.29858456686
Cbr0 netL0 node_ref 2.221486955304943e-08

* Branch 1
Rabr1 node_3 netRa1 23.97092422447678
Lbr1 netRa1 netL1 0.01655505783855915
Rbbr1 netL1 node_ref 24314.77955789861
Cbr1 netL1 node_ref 3.998093983020541e-08

* Branch 2
Rabr2 node_3 netRa2 -80.53191078383787
Lbr2 netRa2 netL2 0.0430884063243866
Rbbr2 netL2 node_ref -28481.82621995759
Cbr2 netL2 node_ref 1.514039473324074e-08

* Branch 3
Rabr3 node_3 netRa3 284.7911106620841
Lbr3 netRa3 netL3 0.03451797738671303
Rbbr3 netL3 node_ref 266153.1416134351
Cbr3 netL3 node_ref 2.463498888694679e-09

* Branch 4
Rabr4 node_3 netRa4 51.35181677247574
Lbr4 netRa4 netL4 0.01661824993789196
Rbbr4 netL4 node_ref 98263.51501565707
Cbr4 netL4 node_ref 4.404482496919189e-09

* Branch 5
Rabr5 node_3 netRa5 -133.93483142158516
Lbr5 netRa5 netL5 0.04242291674017906
Rbbr5 netL5 node_ref -149592.78834168628
Cbr5 netL5 node_ref 1.7061983924393958e-09

* Branch 6
Rabr6 node_3 netRa6 476.9334390075544
Lbr6 netRa6 netL6 0.033604610711336136
Rbbr6 netL6 node_ref 359310.375907067
Cbr6 netL6 node_ref 8.924682559742155e-10

* Branch 7
Rabr7 node_3 netRa7 110.96724584478416
Lbr7 netRa7 netL7 0.01580631360411644
Rbbr7 netL7 node_ref 102498.09162027646
Cbr7 netL7 node_ref 1.662917287657302e-09

* Branch 8
Rabr8 node_3 netRa8 -596.6858836538272
Lbr8 netRa8 netL8 0.04729977250099182
Rbbr8 netL8 node_ref -134389.70192382723
Cbr8 netL8 node_ref 5.48686756683558e-10

* Branch 9
Rabr9 node_3 netRa9 577.5568832916686
Lbr9 netRa9 netL9 0.03249189257621765
Rbbr9 netL9 node_ref 855330.5591527633
Cbr9 netL9 node_ref 4.6460874302326943e-10

* Branch 10
Rabr10 node_3 netRa10 61.07271315221466
Lbr10 netRa10 netL10 0.015984030440449715
Rbbr10 netL10 node_ref 507457.2168351258
Cbr10 netL10 node_ref 8.389822207433891e-10

* Branch 11
Rabr11 node_3 netRa11 111.29626450858697
Lbr11 netRa11 netL11 0.04468223825097084
Rbbr11 netL11 node_ref 2499265.822551149
Cbr11 netL11 node_ref 2.97449223919291e-10

* Branch 12
Rabr12 node_3 netRa12 609.246825849404
Lbr12 netRa12 netL12 0.031282681971788406
Rbbr12 netL12 node_ref 61028624.02375445
Cbr12 netL12 node_ref 2.8909752985160475e-10

* Branch 13
Rabr13 node_3 netRa13 103.61963736973688
Lbr13 netRa13 netL13 0.01568642258644104
Rbbr13 netL13 node_ref 406239.2500308092
Cbr13 netL13 node_ref 5.167552336953745e-10

* Branch 14
Rabr14 node_3 netRa14 51.50012020780365
Lbr14 netRa14 netL14 0.04599593207240105
Rbbr14 netL14 node_ref -40290937.88077229
Cbr14 netL14 node_ref 1.747381220613374e-10

* Branch 15
Rabr15 node_3 netRa15 466.09937405983766
Lbr15 netRa15 netL15 0.030966438353061676
Rbbr15 netL15 node_ref -653521.8212227856
Cbr15 netL15 node_ref 1.940565573658753e-10

* Branch 16
Rabr16 node_3 netRa16 36.20229772498286
Lbr16 netRa16 netL16 0.015594634227454662
Rbbr16 netL16 node_ref 19957307.02570276
Cbr16 netL16 node_ref 3.4782298578574673e-10

* Branch 17
Rabr17 node_3 netRa17 802.21013722832
Lbr17 netRa17 netL17 0.04518767446279526
Rbbr17 netL17 node_ref 514865.8899008287
Cbr17 netL17 node_ref 1.1883822778727674e-10

* Branch 18
Rabr18 node_3 netRa18 -772.8739795137145
Lbr18 netRa18 netL18 0.03216779604554176
Rbbr18 netL18 node_ref -152609.6954652635
Cbr18 netL18 node_ref 1.3192331402624544e-10

* Branch 19
Rabr19 node_3 netRa19 -106.60960160781026
Lbr19 netRa19 netL19 0.015438985079526901
Rbbr19 netL19 node_ref -422236.21560827084
Cbr19 netL19 node_ref 2.5131929904167295e-10

* Branch 20
Rabr20 node_3 netRa20 1910.1162684640065
Lbr20 netRa20 netL20 0.04415206238627434
Rbbr20 netL20 node_ref 277026.0023609452
Cbr20 netL20 node_ref 8.659131497775039e-11

* Branch 21
Rabr21 node_3 netRa21 -6414.511672807723
Lbr21 netRa21 netL21 0.03976304829120636
Rbbr21 netL21 node_ref -73293.8166760016
Cbr21 netL21 node_ref 7.289610629705023e-11

* Branch 22
Rabr22 node_3 netRa22 -321.9703869967046
Lbr22 netRa22 netL22 0.015935653820633888
Rbbr22 netL22 node_ref -238240.7991738014
Cbr22 netL22 node_ref 1.8259449141475423e-10

* Branch 23
Rabr23 node_3 netRa23 1659.6221779954433
Lbr23 netRa23 netL23 0.04173152521252632
Rbbr23 netL23 node_ref 381421.1098806523
Cbr23 netL23 node_ref 6.89703224296523e-11

* Branch 24
Rabr24 node_3 netRa24 572.7548833898331
Lbr24 netRa24 netL24 0.0010093661257997155
Rbbr24 netL24 node_ref 2018.6334125094236
Cbr24 netL24 node_ref 1.2626807262004068e-09

.ends


.end
